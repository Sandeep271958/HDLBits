module top_module(
    input clk,
    input in,
    input areset,
    output out); //
    
    parameter A = 2'b00, B = 2'b01, C = 2'b10, D = 2'b11;
    reg [1:0] state, next_state;
   
    // State transition logic
    always@(*)
        begin
            case(state)
                A: begin 
                    next_state = in ? B : A;
                    out = 0;
                end
                B: begin 
                    next_state = in ? B : C;
                    out = 0;
                end
                C: begin
                    next_state = in ? D : A;
                    out = 0;
                end
                D: begin
                    next_state = in ? B : C;
                    out = 1;
                end
                default: begin
                    next_state = A;
                    out = 0;
                end

            endcase
        end
    
    
    // State flip-flops with asynchronous reset

    always@(posedge clk or posedge areset)
        begin
            if(areset)
                state <= A;
            else
                begin
                   state <= next_state;
                end
            
        end

    // Output logic

endmodule
